CircuitMaker Text
5.6
Probes: 3
R1_2
Transient Analysis
0 404 218 65280
R2_2
Transient Analysis
1 544 217 65535
R3_2
Transient Analysis
2 683 214 16776960
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 10
181 80 1364 405
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 2 0.500000 0.500000
349 176 1532 509
9961490 0
0
6 Title:
5 Name:
0
0
0
20
7 Ground~
168 174 395 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4299 0 0
2
45139.5 0
0
10 Polar Cap~
219 939 165 0 2 5
0 8 4
0
0 0 848 270
3 1uF
10 4 31 12
2 C1
14 -6 28 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
9672 0 0
2
45139.5 0
0
9 Inductor~
219 834 97 0 2 5
0 10 9
0
0 0 848 0
5 0.5mH
-18 -17 17 -9
2 L4
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 0 0 0 0
1 L
7876 0 0
2
45139.5 0
0
6 Diode~
219 687 269 0 2 5
0 3 6
0
0 0 848 90
6 1N3064
12 0 54 8
2 D6
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
6369 0 0
2
45139.5 0
0
6 Diode~
219 682 140 0 2 5
0 6 10
0
0 0 848 90
6 1N3064
12 0 54 8
2 D5
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
9172 0 0
2
45139.5 0
0
6 Diode~
219 548 265 0 2 5
0 4 5
0
0 0 848 90
6 1N3064
12 0 54 8
2 D4
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
7100 0 0
2
45139.5 0
0
6 Diode~
219 543 140 0 2 5
0 5 10
0
0 0 848 90
6 1N3064
12 0 54 8
2 D3
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
3820 0 0
2
45139.5 0
0
6 Diode~
219 402 260 0 2 5
0 4 7
0
0 0 848 90
6 1N3064
12 0 54 8
2 D2
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
7678 0 0
2
45139.5 0
0
6 Diode~
219 400 136 0 2 5
0 7 10
0
0 0 848 90
6 1N3064
12 0 54 8
2 D1
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
961 0 0
2
45139.5 0
0
9 Inductor~
219 152 131 0 2 5
0 11 14
0
0 0 848 0
5 0.1mH
-18 -17 17 -9
2 L3
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 0 0 0 0
1 L
3178 0 0
2
45139.5 0
0
9 Inductor~
219 151 91 0 2 5
0 12 15
0
0 0 848 0
5 0.1mH
-18 -17 17 -9
2 L2
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 0 0 0 0
1 L
3409 0 0
2
45139.5 0
0
9 Inductor~
219 149 55 0 2 5
0 13 16
0
0 0 848 0
5 0.1mH
-18 -17 17 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 0 0 0 0
1 L
3951 0 0
2
45139.5 0
0
11 Signal Gen~
195 258 290 0 64 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1012557331 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 0 250 0.01333 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 250 50 13.33m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8885 0 0
2
45139.5 0
0
11 Signal Gen~
195 175 290 0 64 64
0 12 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1004170870 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 0 250 0.006666 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 250 50 6.666m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3780 0 0
2
45139.5 0
0
11 Signal Gen~
195 87 288 0 19 64
0 13 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
20
1 50 0 250 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 250 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9265 0 0
2
45139.5 0
0
9 Resistor~
219 1053 212 0 2 5
0 4 8
0
0 0 880 90
4 16.5
2 0 30 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9442 0 0
2
45139.5 0
0
9 Resistor~
219 915 97 0 2 5
0 9 8
0
0 0 880 0
2 2m
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9424 0 0
2
45139.5 0
0
9 Resistor~
219 246 132 0 2 5
0 14 6
0
0 0 880 0
2 1m
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9968 0 0
2
45139.5 0
0
9 Resistor~
219 243 87 0 2 5
0 15 5
0
0 0 880 0
2 1m
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9281 0 0
2
45139.5 0
0
9 Resistor~
219 238 52 0 2 5
0 16 7
0
0 0 880 0
2 1m
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8464 0 0
2
45139.5 0
0
26
1 0 3 0 0 4096 0 4 0 0 2 2
687 279
687 285
1 0 3 0 0 8320 0 4 0 0 0 3
687 279
687 295
548 295
1 0 4 0 0 4096 0 6 0 0 11 2
548 275
548 291
2 0 5 0 0 4224 0 19 0 0 19 4
261 87
522 87
522 153
543 153
2 0 6 0 0 12416 0 18 0 0 18 4
264 132
371 132
371 157
682 157
2 1 7 0 0 4224 0 20 9 0 0 4
256 52
390 52
390 146
400 146
2 1 2 0 0 8320 0 13 1 0 0 3
289 295
289 389
174 389
2 1 2 0 0 0 0 14 1 0 0 4
206 295
206 338
174 338
174 389
2 1 2 0 0 0 0 15 1 0 0 4
118 293
139 293
139 389
174 389
2 0 4 0 0 8192 0 2 0 0 11 3
938 172
938 249
1053 249
1 1 4 0 0 8320 0 8 16 0 0 4
402 270
402 291
1053 291
1053 230
2 2 8 0 0 4224 0 17 16 0 0 3
933 97
1053 97
1053 194
2 1 8 0 0 0 0 17 2 0 0 3
933 97
933 155
938 155
2 1 9 0 0 4224 0 3 17 0 0 2
852 97
897 97
2 0 10 0 0 4096 0 5 0 0 17 2
682 130
682 97
2 0 10 0 0 0 0 7 0 0 17 2
543 130
543 97
2 1 10 0 0 8320 0 9 3 0 0 3
400 126
400 97
816 97
1 2 6 0 0 0 0 5 4 0 0 3
682 150
682 259
687 259
1 2 5 0 0 0 0 7 6 0 0 3
543 150
543 255
548 255
1 2 7 0 0 128 0 9 8 0 0 3
400 146
402 146
402 250
1 1 11 0 0 12416 0 10 13 0 0 5
134 131
128 131
128 148
289 148
289 285
1 1 12 0 0 16512 0 11 14 0 0 5
133 91
125 91
125 162
206 162
206 285
1 1 13 0 0 4224 0 15 12 0 0 3
118 283
118 55
131 55
2 1 14 0 0 8320 0 10 18 0 0 3
170 131
170 132
228 132
2 1 15 0 0 4224 0 11 19 0 0 4
169 91
220 91
220 87
225 87
1 2 16 0 0 8320 0 20 12 0 0 3
220 52
220 55
167 55
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
6685644 1079360 100 100 0 0
77 66 977 186
0 74 161 144
977 66
77 66
977 66
977 186
0 0
5.2221e-315 0 5.59737e-315 1.62074e-314 5.2221e-315 5.63882e-315
12385 0
4 0.01 10000
0
6685668 8550976 100 100 0 0
77 66 977 246
0 406 1024 738
977 66
77 66
977 66
977 180
0 0
5.10978e-315 5.02812e-315 5.60223e-315 1.61326e-314 5.10896e-315 5.10896e-315
12409 0
2 0.01 100
4
764 118
0 4 0 0 1	0 27 0 0
356 156
0 7 0 0 3	0 27 0 0
443 153
0 6 0 0 1	0 27 0 0
542 152
0 5 0 0 1	0 27 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
